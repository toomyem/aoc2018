module day04

import utils

fn prepare(input []string) ![]string {
	return input
}

fn solve1(input []string) !string {
	return '1'
}

fn solve2(input []string) !string {
	return '2'
}

pub fn main() ! {
	utils.print_solution(4, prepare, solve1, solve2)!
}
