module main

import day01

pub fn main() {
	day01.main()
}
